// Quick blinking a LED

/* module */
module blinking (

    input CLOCK_50,
    output [7:0] LEDG
    // output LEDG
);

    /* reg */
    // reg data1 = 1'b1;
    reg [32:0] counter;
    reg [7:0] state;
    
    /* assign */
    assign LEDG = state;
    // assign LEDG[1] = data1;
    
    /* always */
    always @ (posedge CLOCK_50) begin
        counter <= counter + 1;
        state <= counter[29:22]; // <------ data to change
    end

endmodule

